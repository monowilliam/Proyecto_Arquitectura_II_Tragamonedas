library verilog;
use verilog.vl_types.all;
entity Mux12_vlg_vec_tst is
end Mux12_vlg_vec_tst;
