library verilog;
use verilog.vl_types.all;
entity Mux14_vlg_vec_tst is
end Mux14_vlg_vec_tst;
