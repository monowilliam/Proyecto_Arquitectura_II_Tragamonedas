library verilog;
use verilog.vl_types.all;
entity memoriaram_vlg_vec_tst is
end memoriaram_vlg_vec_tst;
