library verilog;
use verilog.vl_types.all;
entity Registro_vlg_vec_tst is
end Registro_vlg_vec_tst;
