library verilog;
use verilog.vl_types.all;
entity sieteS_vlg_vec_tst is
end sieteS_vlg_vec_tst;
