library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity memoria is generic(
	BusInstruc: natural);
port(
	clk : in std_logic;
	address: in integer range 0 to 255;
	data_out : out std_logic_vector(BusInstruc-1 downto 0)
);
end entity;

architecture mem_arc of memoria is
signal reg_address: integer range 0 to 255;
type memoria is array(0 to 255) of std_logic_vector(BusInstruc-1 downto 0);
signal my_rom : memoria   := (
	0 => "00010100000000000000000000",
	1 => "00010111000000000000000000", 
	2 => "00000111000000000000000000", 
	3 => "01010111011100000000000000", 
	4 => "01100111000000000000000000",
--	5 => "00010100011100000000000000",
--	6 => "00010111000000000000000001",
--	7 => "00000111000000000000000000",
--	8 => "01010111011100000000000000",
--	9 => "10000111010000000000000110",
--	10 => "01100111000000000000000110",
--	11 => "01000111000000000000000001",
--	12 => "00010101011100000000000000",
--	13 => "00011000000000000000000001",
--	14 => "10010100010100000000000000",
--	15 => "01000100000000000000000000",
--	16 => "00010111000000000000000011",
--	17 => "11000111000000000000000000",
--	18 => "00010110000000000000000001",
--	19 => "01000110000000000000000010",
--	20 => "01010111011100000000000000",
--	21 => "01110111000000000000011010",
--	22 => "00011000000000000000000000",
--	23 => "10111000000000000000000000",
--	24 => "01110100000000000000000110",
--	25 => "10100000000000000000000000",
--	26 => "00110110001100000000000000",
--	27 => "01000110000000000000000010",
--	28 => "00110101011000000000000000",
--	29 => "00100100010100000000000000",
--	30 => "00011000000000000000000000",
--	31 => "10111000000000000000000000",
--	32 => "01000100000000000000000000",
--	33 => "01000000000000000000000001",
--	34 => "10100000000000000000000110",
	others => "11111111111111111111111111"
);	
begin
	process(clk) is
	begin
		if(rising_edge(clk)) then
			reg_address <= address;
		end if;
	end process;
	data_out <= my_rom(reg_address);
end architecture;