library verilog;
use verilog.vl_types.all;
entity sumPC_vlg_vec_tst is
end sumPC_vlg_vec_tst;
