library verilog;
use verilog.vl_types.all;
entity UC_vlg_vec_tst is
end UC_vlg_vec_tst;
