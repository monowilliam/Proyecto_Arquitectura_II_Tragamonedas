library verilog;
use verilog.vl_types.all;
entity mostrar_vlg_vec_tst is
end mostrar_vlg_vec_tst;
