library verilog;
use verilog.vl_types.all;
entity PCounter_vlg_vec_tst is
end PCounter_vlg_vec_tst;
