library verilog;
use verilog.vl_types.all;
entity randomSegmento_vlg_vec_tst is
end randomSegmento_vlg_vec_tst;
