library verilog;
use verilog.vl_types.all;
entity Principal_vlg_vec_tst is
end Principal_vlg_vec_tst;
